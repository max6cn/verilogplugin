// this is a comment
module aaabb ;
endmodule
// this is a test
module abc;
endmodule

// this is a test
module abc;
endmmodule

module a;
endmodule
